library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sigmoid_lut_2048 is
  port (
    address : in  std_logic_vector(10 downto 0);
    dds_out : out std_logic_vector(15 downto 0) 
  );
end sigmoid_lut_2048;


-- Output between [-11; +11], rapresented with fixed point
-- Need for 1 bit for integer, last 15 bit for float rapresentation
-- Reach the LSB method
-- 
-- LSB(in) = (11)/(2^11 - 1) = 0.00537371763556424035173424523693
-- LSB(out) = (1)/(2^15 - 1) = 3.0518509475997192297128208258309e-5
-- inputs -> [-11, +11] 
-- outputs -> [0, 1]
-- Q(f(x)) = round(f(x)/LSB(out))*LSB(out)
-- 
--
-- What to store in the lut? round(f(x)/LSB(out)) for x in [0; 2047]*LSB(in)

architecture rtl of sigmoid_lut_2048 is
type LUT_t is array (natural range 0 to 2047) of integer;
constant LUT: LUT_t := (
    0 => 16384,
    1 => 16512,
    2 => 16640,
    3 => 16768,
    4 => 16896,
    5 => 17023,
    6 => 17151,
    7 => 17279,
    8 => 17407,
    9 => 17534,
    10 => 17661,
    11 => 17789,
    12 => 17916,
    13 => 18043,
    14 => 18169,
    15 => 18296,
    16 => 18422,
    17 => 18548,
    18 => 18673,
    19 => 18799,
    20 => 18924,
    21 => 19049,
    22 => 19173,
    23 => 19298,
    24 => 19421,
    25 => 19545,
    26 => 19668,
    27 => 19791,
    28 => 19913,
    29 => 20035,
    30 => 20156,
    31 => 20277,
    32 => 20398,
    33 => 20518,
    34 => 20638,
    35 => 20757,
    36 => 20876,
    37 => 20994,
    38 => 21112,
    39 => 21229,
    40 => 21345,
    41 => 21461,
    42 => 21577,
    43 => 21692,
    44 => 21806,
    45 => 21920,
    46 => 22033,
    47 => 22145,
    48 => 22257,
    49 => 22369,
    50 => 22479,
    51 => 22589,
    52 => 22699,
    53 => 22807,
    54 => 22915,
    55 => 23023,
    56 => 23129,
    57 => 23235,
    58 => 23341,
    59 => 23445,
    60 => 23549,
    61 => 23652,
    62 => 23755,
    63 => 23857,
    64 => 23958,
    65 => 24058,
    66 => 24158,
    67 => 24257,
    68 => 24355,
    69 => 24452,
    70 => 24549,
    71 => 24645,
    72 => 24740,
    73 => 24834,
    74 => 24928,
    75 => 25020,
    76 => 25113,
    77 => 25204,
    78 => 25294,
    79 => 25384,
    80 => 25473,
    81 => 25562,
    82 => 25649,
    83 => 25736,
    84 => 25822,
    85 => 25907,
    86 => 25991,
    87 => 26075,
    88 => 26158,
    89 => 26240,
    90 => 26321,
    91 => 26402,
    92 => 26482,
    93 => 26561,
    94 => 26639,
    95 => 26716,
    96 => 26793,
    97 => 26869,
    98 => 26944,
    99 => 27019,
    100 => 27092,
    101 => 27165,
    102 => 27238,
    103 => 27309,
    104 => 27380,
    105 => 27450,
    106 => 27519,
    107 => 27588,
    108 => 27655,
    109 => 27723,
    110 => 27789,
    111 => 27855,
    112 => 27919,
    113 => 27984,
    114 => 28047,
    115 => 28110,
    116 => 28172,
    117 => 28234,
    118 => 28294,
    119 => 28354,
    120 => 28414,
    121 => 28472,
    122 => 28530,
    123 => 28588,
    124 => 28644,
    125 => 28700,
    126 => 28756,
    127 => 28810,
    128 => 28864,
    129 => 28918,
    130 => 28971,
    131 => 29023,
    132 => 29074,
    133 => 29125,
    134 => 29176,
    135 => 29225,
    136 => 29274,
    137 => 29323,
    138 => 29371,
    139 => 29418,
    140 => 29465,
    141 => 29511,
    142 => 29556,
    143 => 29601,
    144 => 29646,
    145 => 29690,
    146 => 29733,
    147 => 29776,
    148 => 29818,
    149 => 29860,
    150 => 29901,
    151 => 29941,
    152 => 29982,
    153 => 30021,
    154 => 30060,
    155 => 30099,
    156 => 30137,
    157 => 30174,
    158 => 30211,
    159 => 30248,
    160 => 30284,
    161 => 30320,
    162 => 30355,
    163 => 30390,
    164 => 30424,
    165 => 30458,
    166 => 30491,
    167 => 30524,
    168 => 30556,
    169 => 30588,
    170 => 30620,
    171 => 30651,
    172 => 30682,
    173 => 30712,
    174 => 30742,
    175 => 30772,
    176 => 30801,
    177 => 30829,
    178 => 30858,
    179 => 30886,
    180 => 30913,
    181 => 30940,
    182 => 30967,
    183 => 30993,
    184 => 31019,
    185 => 31045,
    186 => 31070,
    187 => 31095,
    188 => 31120,
    189 => 31144,
    190 => 31168,
    191 => 31192,
    192 => 31215,
    193 => 31238,
    194 => 31261,
    195 => 31283,
    196 => 31305,
    197 => 31327,
    198 => 31348,
    199 => 31369,
    200 => 31390,
    201 => 31410,
    202 => 31431,
    203 => 31450,
    204 => 31470,
    205 => 31489,
    206 => 31508,
    207 => 31527,
    208 => 31546,
    209 => 31564,
    210 => 31582,
    211 => 31600,
    212 => 31617,
    213 => 31634,
    214 => 31651,
    215 => 31668,
    216 => 31685,
    217 => 31701,
    218 => 31717,
    219 => 31733,
    220 => 31748,
    221 => 31763,
    222 => 31779,
    223 => 31793,
    224 => 31808,
    225 => 31823,
    226 => 31837,
    227 => 31851,
    228 => 31865,
    229 => 31878,
    230 => 31892,
    231 => 31905,
    232 => 31918,
    233 => 31931,
    234 => 31943,
    235 => 31956,
    236 => 31968,
    237 => 31980,
    238 => 31992,
    239 => 32004,
    240 => 32015,
    241 => 32027,
    242 => 32038,
    243 => 32049,
    244 => 32060,
    245 => 32071,
    246 => 32081,
    247 => 32092,
    248 => 32102,
    249 => 32112,
    250 => 32122,
    251 => 32132,
    252 => 32142,
    253 => 32151,
    254 => 32160,
    255 => 32170,
    256 => 32179,
    257 => 32188,
    258 => 32197,
    259 => 32205,
    260 => 32214,
    261 => 32222,
    262 => 32231,
    263 => 32239,
    264 => 32247,
    265 => 32255,
    266 => 32263,
    267 => 32270,
    268 => 32278,
    269 => 32285,
    270 => 32293,
    271 => 32300,
    272 => 32307,
    273 => 32314,
    274 => 32321,
    275 => 32328,
    276 => 32335,
    277 => 32341,
    278 => 32348,
    279 => 32354,
    280 => 32361,
    281 => 32367,
    282 => 32373,
    283 => 32379,
    284 => 32385,
    285 => 32391,
    286 => 32396,
    287 => 32402,
    288 => 32408,
    289 => 32413,
    290 => 32419,
    291 => 32424,
    292 => 32429,
    293 => 32435,
    294 => 32440,
    295 => 32445,
    296 => 32450,
    297 => 32454,
    298 => 32459,
    299 => 32464,
    300 => 32469,
    301 => 32473,
    302 => 32478,
    303 => 32482,
    304 => 32487,
    305 => 32491,
    306 => 32495,
    307 => 32499,
    308 => 32503,
    309 => 32508,
    310 => 32511,
    311 => 32515,
    312 => 32519,
    313 => 32523,
    314 => 32527,
    315 => 32531,
    316 => 32534,
    317 => 32538,
    318 => 32541,
    319 => 32545,
    320 => 32548,
    321 => 32552,
    322 => 32555,
    323 => 32558,
    324 => 32561,
    325 => 32565,
    326 => 32568,
    327 => 32571,
    328 => 32574,
    329 => 32577,
    330 => 32580,
    331 => 32583,
    332 => 32585,
    333 => 32588,
    334 => 32591,
    335 => 32594,
    336 => 32596,
    337 => 32599,
    338 => 32602,
    339 => 32604,
    340 => 32607,
    341 => 32609,
    342 => 32612,
    343 => 32614,
    344 => 32616,
    345 => 32619,
    346 => 32621,
    347 => 32623,
    348 => 32625,
    349 => 32628,
    350 => 32630,
    351 => 32632,
    352 => 32634,
    353 => 32636,
    354 => 32638,
    355 => 32640,
    356 => 32642,
    357 => 32644,
    358 => 32646,
    359 => 32648,
    360 => 32650,
    361 => 32651,
    362 => 32653,
    363 => 32655,
    364 => 32657,
    365 => 32658,
    366 => 32660,
    367 => 32662,
    368 => 32663,
    369 => 32665,
    370 => 32667,
    371 => 32668,
    372 => 32670,
    373 => 32671,
    374 => 32673,
    375 => 32674,
    376 => 32675,
    377 => 32677,
    378 => 32678,
    379 => 32680,
    380 => 32681,
    381 => 32682,
    382 => 32684,
    383 => 32685,
    384 => 32686,
    385 => 32687,
    386 => 32689,
    387 => 32690,
    388 => 32691,
    389 => 32692,
    390 => 32693,
    391 => 32695,
    392 => 32696,
    393 => 32697,
    394 => 32698,
    395 => 32699,
    396 => 32700,
    397 => 32701,
    398 => 32702,
    399 => 32703,
    400 => 32704,
    401 => 32705,
    402 => 32706,
    403 => 32707,
    404 => 32708,
    405 => 32709,
    406 => 32710,
    407 => 32711,
    408 => 32711,
    409 => 32712,
    410 => 32713,
    411 => 32714,
    412 => 32715,
    413 => 32716,
    414 => 32716,
    415 => 32717,
    416 => 32718,
    417 => 32719,
    418 => 32719,
    419 => 32720,
    420 => 32721,
    421 => 32722,
    422 => 32722,
    423 => 32723,
    424 => 32724,
    425 => 32724,
    426 => 32725,
    427 => 32726,
    428 => 32726,
    429 => 32727,
    430 => 32728,
    431 => 32728,
    432 => 32729,
    433 => 32729,
    434 => 32730,
    435 => 32731,
    436 => 32731,
    437 => 32732,
    438 => 32732,
    439 => 32733,
    440 => 32733,
    441 => 32734,
    442 => 32734,
    443 => 32735,
    444 => 32735,
    445 => 32736,
    446 => 32736,
    447 => 32737,
    448 => 32737,
    449 => 32738,
    450 => 32738,
    451 => 32739,
    452 => 32739,
    453 => 32739,
    454 => 32740,
    455 => 32740,
    456 => 32741,
    457 => 32741,
    458 => 32742,
    459 => 32742,
    460 => 32742,
    461 => 32743,
    462 => 32743,
    463 => 32743,
    464 => 32744,
    465 => 32744,
    466 => 32745,
    467 => 32745,
    468 => 32745,
    469 => 32746,
    470 => 32746,
    471 => 32746,
    472 => 32747,
    473 => 32747,
    474 => 32747,
    475 => 32747,
    476 => 32748,
    477 => 32748,
    478 => 32748,
    479 => 32749,
    480 => 32749,
    481 => 32749,
    482 => 32750,
    483 => 32750,
    484 => 32750,
    485 => 32750,
    486 => 32751,
    487 => 32751,
    488 => 32751,
    489 => 32751,
    490 => 32752,
    491 => 32752,
    492 => 32752,
    493 => 32752,
    494 => 32752,
    495 => 32753,
    496 => 32753,
    497 => 32753,
    498 => 32753,
    499 => 32754,
    500 => 32754,
    501 => 32754,
    502 => 32754,
    503 => 32754,
    504 => 32755,
    505 => 32755,
    506 => 32755,
    507 => 32755,
    508 => 32755,
    509 => 32756,
    510 => 32756,
    511 => 32756,
    512 => 32756,
    513 => 32756,
    514 => 32756,
    515 => 32757,
    516 => 32757,
    517 => 32757,
    518 => 32757,
    519 => 32757,
    520 => 32757,
    521 => 32757,
    522 => 32758,
    523 => 32758,
    524 => 32758,
    525 => 32758,
    526 => 32758,
    527 => 32758,
    528 => 32758,
    529 => 32759,
    530 => 32759,
    531 => 32759,
    532 => 32759,
    533 => 32759,
    534 => 32759,
    535 => 32759,
    536 => 32759,
    537 => 32760,
    538 => 32760,
    539 => 32760,
    540 => 32760,
    541 => 32760,
    542 => 32760,
    543 => 32760,
    544 => 32760,
    545 => 32760,
    546 => 32761,
    547 => 32761,
    548 => 32761,
    549 => 32761,
    550 => 32761,
    551 => 32761,
    552 => 32761,
    553 => 32761,
    554 => 32761,
    555 => 32761,
    556 => 32761,
    557 => 32762,
    558 => 32762,
    559 => 32762,
    560 => 32762,
    561 => 32762,
    562 => 32762,
    563 => 32762,
    564 => 32762,
    565 => 32762,
    566 => 32762,
    567 => 32762,
    568 => 32762,
    569 => 32763,
    570 => 32763,
    571 => 32763,
    572 => 32763,
    573 => 32763,
    574 => 32763,
    575 => 32763,
    576 => 32763,
    577 => 32763,
    578 => 32763,
    579 => 32763,
    580 => 32763,
    581 => 32763,
    582 => 32763,
    583 => 32763,
    584 => 32763,
    585 => 32764,
    586 => 32764,
    587 => 32764,
    588 => 32764,
    589 => 32764,
    590 => 32764,
    591 => 32764,
    592 => 32764,
    593 => 32764,
    594 => 32764,
    595 => 32764,
    596 => 32764,
    597 => 32764,
    598 => 32764,
    599 => 32764,
    600 => 32764,
    601 => 32764,
    602 => 32764,
    603 => 32764,
    604 => 32764,
    605 => 32764,
    606 => 32764,
    607 => 32765,
    608 => 32765,
    609 => 32765,
    610 => 32765,
    611 => 32765,
    612 => 32765,
    613 => 32765,
    614 => 32765,
    615 => 32765,
    616 => 32765,
    617 => 32765,
    618 => 32765,
    619 => 32765,
    620 => 32765,
    621 => 32765,
    622 => 32765,
    623 => 32765,
    624 => 32765,
    625 => 32765,
    626 => 32765,
    627 => 32765,
    628 => 32765,
    629 => 32765,
    630 => 32765,
    631 => 32765,
    632 => 32765,
    633 => 32765,
    634 => 32765,
    635 => 32765,
    636 => 32765,
    637 => 32765,
    638 => 32765,
    639 => 32765,
    640 => 32766,
    641 => 32766,
    642 => 32766,
    643 => 32766,
    644 => 32766,
    645 => 32766,
    646 => 32766,
    647 => 32766,
    648 => 32766,
    649 => 32766,
    650 => 32766,
    651 => 32766,
    652 => 32766,
    653 => 32766,
    654 => 32766,
    655 => 32766,
    656 => 32766,
    657 => 32766,
    658 => 32766,
    659 => 32766,
    660 => 32766,
    661 => 32766,
    662 => 32766,
    663 => 32766,
    664 => 32766,
    665 => 32766,
    666 => 32766,
    667 => 32766,
    668 => 32766,
    669 => 32766,
    670 => 32766,
    671 => 32766,
    672 => 32766,
    673 => 32766,
    674 => 32766,
    675 => 32766,
    676 => 32766,
    677 => 32766,
    678 => 32766,
    679 => 32766,
    680 => 32766,
    681 => 32766,
    682 => 32766,
    683 => 32766,
    684 => 32766,
    685 => 32766,
    686 => 32766,
    687 => 32766,
    688 => 32766,
    689 => 32766,
    690 => 32766,
    691 => 32766,
    692 => 32766,
    693 => 32766,
    694 => 32766,
    695 => 32766,
    696 => 32766,
    697 => 32766,
    698 => 32766,
    699 => 32766,
    700 => 32766,
    701 => 32766,
    702 => 32766,
    703 => 32766,
    704 => 32766,
    705 => 32766,
    706 => 32766,
    707 => 32766,
    708 => 32766,
    709 => 32766,
    710 => 32767,
    711 => 32767,
    712 => 32767,
    713 => 32767,
    714 => 32767,
    715 => 32767,
    716 => 32767,
    717 => 32767,
    718 => 32767,
    719 => 32767,
    720 => 32767,
    721 => 32767,
    722 => 32767,
    723 => 32767,
    724 => 32767,
    725 => 32767,
    726 => 32767,
    727 => 32767,
    728 => 32767,
    729 => 32767,
    730 => 32767,
    731 => 32767,
    732 => 32767,
    733 => 32767,
    734 => 32767,
    735 => 32767,
    736 => 32767,
    737 => 32767,
    738 => 32767,
    739 => 32767,
    740 => 32767,
    741 => 32767,
    742 => 32767,
    743 => 32767,
    744 => 32767,
    745 => 32767,
    746 => 32767,
    747 => 32767,
    748 => 32767,
    749 => 32767,
    750 => 32767,
    751 => 32767,
    752 => 32767,
    753 => 32767,
    754 => 32767,
    755 => 32767,
    756 => 32767,
    757 => 32767,
    758 => 32767,
    759 => 32767,
    760 => 32767,
    761 => 32767,
    762 => 32767,
    763 => 32767,
    764 => 32767,
    765 => 32767,
    766 => 32767,
    767 => 32767,
    768 => 32767,
    769 => 32767,
    770 => 32767,
    771 => 32767,
    772 => 32767,
    773 => 32767,
    774 => 32767,
    775 => 32767,
    776 => 32767,
    777 => 32767,
    778 => 32767,
    779 => 32767,
    780 => 32767,
    781 => 32767,
    782 => 32767,
    783 => 32767,
    784 => 32767,
    785 => 32767,
    786 => 32767,
    787 => 32767,
    788 => 32767,
    789 => 32767,
    790 => 32767,
    791 => 32767,
    792 => 32767,
    793 => 32767,
    794 => 32767,
    795 => 32767,
    796 => 32767,
    797 => 32767,
    798 => 32767,
    799 => 32767,
    800 => 32767,
    801 => 32767,
    802 => 32767,
    803 => 32767,
    804 => 32767,
    805 => 32767,
    806 => 32767,
    807 => 32767,
    808 => 32767,
    809 => 32767,
    810 => 32767,
    811 => 32767,
    812 => 32767,
    813 => 32767,
    814 => 32767,
    815 => 32767,
    816 => 32767,
    817 => 32767,
    818 => 32767,
    819 => 32767,
    820 => 32767,
    821 => 32767,
    822 => 32767,
    823 => 32767,
    824 => 32767,
    825 => 32767,
    826 => 32767,
    827 => 32767,
    828 => 32767,
    829 => 32767,
    830 => 32767,
    831 => 32767,
    832 => 32767,
    833 => 32767,
    834 => 32767,
    835 => 32767,
    836 => 32767,
    837 => 32767,
    838 => 32767,
    839 => 32767,
    840 => 32767,
    841 => 32767,
    842 => 32767,
    843 => 32767,
    844 => 32767,
    845 => 32767,
    846 => 32767,
    847 => 32767,
    848 => 32767,
    849 => 32767,
    850 => 32767,
    851 => 32767,
    852 => 32767,
    853 => 32767,
    854 => 32767,
    855 => 32767,
    856 => 32767,
    857 => 32767,
    858 => 32767,
    859 => 32767,
    860 => 32767,
    861 => 32767,
    862 => 32767,
    863 => 32767,
    864 => 32767,
    865 => 32767,
    866 => 32767,
    867 => 32767,
    868 => 32767,
    869 => 32767,
    870 => 32767,
    871 => 32767,
    872 => 32767,
    873 => 32767,
    874 => 32767,
    875 => 32767,
    876 => 32767,
    877 => 32767,
    878 => 32767,
    879 => 32767,
    880 => 32767,
    881 => 32767,
    882 => 32767,
    883 => 32767,
    884 => 32767,
    885 => 32767,
    886 => 32767,
    887 => 32767,
    888 => 32767,
    889 => 32767,
    890 => 32767,
    891 => 32767,
    892 => 32767,
    893 => 32767,
    894 => 32767,
    895 => 32767,
    896 => 32767,
    897 => 32767,
    898 => 32767,
    899 => 32767,
    900 => 32767,
    901 => 32767,
    902 => 32767,
    903 => 32767,
    904 => 32767,
    905 => 32767,
    906 => 32767,
    907 => 32767,
    908 => 32767,
    909 => 32767,
    910 => 32767,
    911 => 32767,
    912 => 32767,
    913 => 32767,
    914 => 32767,
    915 => 32767,
    916 => 32767,
    917 => 32767,
    918 => 32767,
    919 => 32767,
    920 => 32767,
    921 => 32767,
    922 => 32767,
    923 => 32767,
    924 => 32767,
    925 => 32767,
    926 => 32767,
    927 => 32767,
    928 => 32767,
    929 => 32767,
    930 => 32767,
    931 => 32767,
    932 => 32767,
    933 => 32767,
    934 => 32767,
    935 => 32767,
    936 => 32767,
    937 => 32767,
    938 => 32767,
    939 => 32767,
    940 => 32767,
    941 => 32767,
    942 => 32767,
    943 => 32767,
    944 => 32767,
    945 => 32767,
    946 => 32767,
    947 => 32767,
    948 => 32767,
    949 => 32767,
    950 => 32767,
    951 => 32767,
    952 => 32767,
    953 => 32767,
    954 => 32767,
    955 => 32767,
    956 => 32767,
    957 => 32767,
    958 => 32767,
    959 => 32767,
    960 => 32767,
    961 => 32767,
    962 => 32767,
    963 => 32767,
    964 => 32767,
    965 => 32767,
    966 => 32767,
    967 => 32767,
    968 => 32767,
    969 => 32767,
    970 => 32767,
    971 => 32767,
    972 => 32767,
    973 => 32767,
    974 => 32767,
    975 => 32767,
    976 => 32767,
    977 => 32767,
    978 => 32767,
    979 => 32767,
    980 => 32767,
    981 => 32767,
    982 => 32767,
    983 => 32767,
    984 => 32767,
    985 => 32767,
    986 => 32767,
    987 => 32767,
    988 => 32767,
    989 => 32767,
    990 => 32767,
    991 => 32767,
    992 => 32767,
    993 => 32767,
    994 => 32767,
    995 => 32767,
    996 => 32767,
    997 => 32767,
    998 => 32767,
    999 => 32767,
    1000 => 32767,
    1001 => 32767,
    1002 => 32767,
    1003 => 32767,
    1004 => 32767,
    1005 => 32767,
    1006 => 32767,
    1007 => 32767,
    1008 => 32767,
    1009 => 32767,
    1010 => 32767,
    1011 => 32767,
    1012 => 32767,
    1013 => 32767,
    1014 => 32767,
    1015 => 32767,
    1016 => 32767,
    1017 => 32767,
    1018 => 32767,
    1019 => 32767,
    1020 => 32767,
    1021 => 32767,
    1022 => 32767,
    1023 => 32767,
    1024 => 32767,
    1025 => 32767,
    1026 => 32767,
    1027 => 32767,
    1028 => 32767,
    1029 => 32767,
    1030 => 32767,
    1031 => 32767,
    1032 => 32767,
    1033 => 32767,
    1034 => 32767,
    1035 => 32767,
    1036 => 32767,
    1037 => 32767,
    1038 => 32767,
    1039 => 32767,
    1040 => 32767,
    1041 => 32767,
    1042 => 32767,
    1043 => 32767,
    1044 => 32767,
    1045 => 32767,
    1046 => 32767,
    1047 => 32767,
    1048 => 32767,
    1049 => 32767,
    1050 => 32767,
    1051 => 32767,
    1052 => 32767,
    1053 => 32767,
    1054 => 32767,
    1055 => 32767,
    1056 => 32767,
    1057 => 32767,
    1058 => 32767,
    1059 => 32767,
    1060 => 32767,
    1061 => 32767,
    1062 => 32767,
    1063 => 32767,
    1064 => 32767,
    1065 => 32767,
    1066 => 32767,
    1067 => 32767,
    1068 => 32767,
    1069 => 32767,
    1070 => 32767,
    1071 => 32767,
    1072 => 32767,
    1073 => 32767,
    1074 => 32767,
    1075 => 32767,
    1076 => 32767,
    1077 => 32767,
    1078 => 32767,
    1079 => 32767,
    1080 => 32767,
    1081 => 32767,
    1082 => 32767,
    1083 => 32767,
    1084 => 32767,
    1085 => 32767,
    1086 => 32767,
    1087 => 32767,
    1088 => 32767,
    1089 => 32767,
    1090 => 32767,
    1091 => 32767,
    1092 => 32767,
    1093 => 32767,
    1094 => 32767,
    1095 => 32767,
    1096 => 32767,
    1097 => 32767,
    1098 => 32767,
    1099 => 32767,
    1100 => 32767,
    1101 => 32767,
    1102 => 32767,
    1103 => 32767,
    1104 => 32767,
    1105 => 32767,
    1106 => 32767,
    1107 => 32767,
    1108 => 32767,
    1109 => 32767,
    1110 => 32767,
    1111 => 32767,
    1112 => 32767,
    1113 => 32767,
    1114 => 32767,
    1115 => 32767,
    1116 => 32767,
    1117 => 32767,
    1118 => 32767,
    1119 => 32767,
    1120 => 32767,
    1121 => 32767,
    1122 => 32767,
    1123 => 32767,
    1124 => 32767,
    1125 => 32767,
    1126 => 32767,
    1127 => 32767,
    1128 => 32767,
    1129 => 32767,
    1130 => 32767,
    1131 => 32767,
    1132 => 32767,
    1133 => 32767,
    1134 => 32767,
    1135 => 32767,
    1136 => 32767,
    1137 => 32767,
    1138 => 32767,
    1139 => 32767,
    1140 => 32767,
    1141 => 32767,
    1142 => 32767,
    1143 => 32767,
    1144 => 32767,
    1145 => 32767,
    1146 => 32767,
    1147 => 32767,
    1148 => 32767,
    1149 => 32767,
    1150 => 32767,
    1151 => 32767,
    1152 => 32767,
    1153 => 32767,
    1154 => 32767,
    1155 => 32767,
    1156 => 32767,
    1157 => 32767,
    1158 => 32767,
    1159 => 32767,
    1160 => 32767,
    1161 => 32767,
    1162 => 32767,
    1163 => 32767,
    1164 => 32767,
    1165 => 32767,
    1166 => 32767,
    1167 => 32767,
    1168 => 32767,
    1169 => 32767,
    1170 => 32767,
    1171 => 32767,
    1172 => 32767,
    1173 => 32767,
    1174 => 32767,
    1175 => 32767,
    1176 => 32767,
    1177 => 32767,
    1178 => 32767,
    1179 => 32767,
    1180 => 32767,
    1181 => 32767,
    1182 => 32767,
    1183 => 32767,
    1184 => 32767,
    1185 => 32767,
    1186 => 32767,
    1187 => 32767,
    1188 => 32767,
    1189 => 32767,
    1190 => 32767,
    1191 => 32767,
    1192 => 32767,
    1193 => 32767,
    1194 => 32767,
    1195 => 32767,
    1196 => 32767,
    1197 => 32767,
    1198 => 32767,
    1199 => 32767,
    1200 => 32767,
    1201 => 32767,
    1202 => 32767,
    1203 => 32767,
    1204 => 32767,
    1205 => 32767,
    1206 => 32767,
    1207 => 32767,
    1208 => 32767,
    1209 => 32767,
    1210 => 32767,
    1211 => 32767,
    1212 => 32767,
    1213 => 32767,
    1214 => 32767,
    1215 => 32767,
    1216 => 32767,
    1217 => 32767,
    1218 => 32767,
    1219 => 32767,
    1220 => 32767,
    1221 => 32767,
    1222 => 32767,
    1223 => 32767,
    1224 => 32767,
    1225 => 32767,
    1226 => 32767,
    1227 => 32767,
    1228 => 32767,
    1229 => 32767,
    1230 => 32767,
    1231 => 32767,
    1232 => 32767,
    1233 => 32767,
    1234 => 32767,
    1235 => 32767,
    1236 => 32767,
    1237 => 32767,
    1238 => 32767,
    1239 => 32767,
    1240 => 32767,
    1241 => 32767,
    1242 => 32767,
    1243 => 32767,
    1244 => 32767,
    1245 => 32767,
    1246 => 32767,
    1247 => 32767,
    1248 => 32767,
    1249 => 32767,
    1250 => 32767,
    1251 => 32767,
    1252 => 32767,
    1253 => 32767,
    1254 => 32767,
    1255 => 32767,
    1256 => 32767,
    1257 => 32767,
    1258 => 32767,
    1259 => 32767,
    1260 => 32767,
    1261 => 32767,
    1262 => 32767,
    1263 => 32767,
    1264 => 32767,
    1265 => 32767,
    1266 => 32767,
    1267 => 32767,
    1268 => 32767,
    1269 => 32767,
    1270 => 32767,
    1271 => 32767,
    1272 => 32767,
    1273 => 32767,
    1274 => 32767,
    1275 => 32767,
    1276 => 32767,
    1277 => 32767,
    1278 => 32767,
    1279 => 32767,
    1280 => 32767,
    1281 => 32767,
    1282 => 32767,
    1283 => 32767,
    1284 => 32767,
    1285 => 32767,
    1286 => 32767,
    1287 => 32767,
    1288 => 32767,
    1289 => 32767,
    1290 => 32767,
    1291 => 32767,
    1292 => 32767,
    1293 => 32767,
    1294 => 32767,
    1295 => 32767,
    1296 => 32767,
    1297 => 32767,
    1298 => 32767,
    1299 => 32767,
    1300 => 32767,
    1301 => 32767,
    1302 => 32767,
    1303 => 32767,
    1304 => 32767,
    1305 => 32767,
    1306 => 32767,
    1307 => 32767,
    1308 => 32767,
    1309 => 32767,
    1310 => 32767,
    1311 => 32767,
    1312 => 32767,
    1313 => 32767,
    1314 => 32767,
    1315 => 32767,
    1316 => 32767,
    1317 => 32767,
    1318 => 32767,
    1319 => 32767,
    1320 => 32767,
    1321 => 32767,
    1322 => 32767,
    1323 => 32767,
    1324 => 32767,
    1325 => 32767,
    1326 => 32767,
    1327 => 32767,
    1328 => 32767,
    1329 => 32767,
    1330 => 32767,
    1331 => 32767,
    1332 => 32767,
    1333 => 32767,
    1334 => 32767,
    1335 => 32767,
    1336 => 32767,
    1337 => 32767,
    1338 => 32767,
    1339 => 32767,
    1340 => 32767,
    1341 => 32767,
    1342 => 32767,
    1343 => 32767,
    1344 => 32767,
    1345 => 32767,
    1346 => 32767,
    1347 => 32767,
    1348 => 32767,
    1349 => 32767,
    1350 => 32767,
    1351 => 32767,
    1352 => 32767,
    1353 => 32767,
    1354 => 32767,
    1355 => 32767,
    1356 => 32767,
    1357 => 32767,
    1358 => 32767,
    1359 => 32767,
    1360 => 32767,
    1361 => 32767,
    1362 => 32767,
    1363 => 32767,
    1364 => 32767,
    1365 => 32767,
    1366 => 32767,
    1367 => 32767,
    1368 => 32767,
    1369 => 32767,
    1370 => 32767,
    1371 => 32767,
    1372 => 32767,
    1373 => 32767,
    1374 => 32767,
    1375 => 32767,
    1376 => 32767,
    1377 => 32767,
    1378 => 32767,
    1379 => 32767,
    1380 => 32767,
    1381 => 32767,
    1382 => 32767,
    1383 => 32767,
    1384 => 32767,
    1385 => 32767,
    1386 => 32767,
    1387 => 32767,
    1388 => 32767,
    1389 => 32767,
    1390 => 32767,
    1391 => 32767,
    1392 => 32767,
    1393 => 32767,
    1394 => 32767,
    1395 => 32767,
    1396 => 32767,
    1397 => 32767,
    1398 => 32767,
    1399 => 32767,
    1400 => 32767,
    1401 => 32767,
    1402 => 32767,
    1403 => 32767,
    1404 => 32767,
    1405 => 32767,
    1406 => 32767,
    1407 => 32767,
    1408 => 32767,
    1409 => 32767,
    1410 => 32767,
    1411 => 32767,
    1412 => 32767,
    1413 => 32767,
    1414 => 32767,
    1415 => 32767,
    1416 => 32767,
    1417 => 32767,
    1418 => 32767,
    1419 => 32767,
    1420 => 32767,
    1421 => 32767,
    1422 => 32767,
    1423 => 32767,
    1424 => 32767,
    1425 => 32767,
    1426 => 32767,
    1427 => 32767,
    1428 => 32767,
    1429 => 32767,
    1430 => 32767,
    1431 => 32767,
    1432 => 32767,
    1433 => 32767,
    1434 => 32767,
    1435 => 32767,
    1436 => 32767,
    1437 => 32767,
    1438 => 32767,
    1439 => 32767,
    1440 => 32767,
    1441 => 32767,
    1442 => 32767,
    1443 => 32767,
    1444 => 32767,
    1445 => 32767,
    1446 => 32767,
    1447 => 32767,
    1448 => 32767,
    1449 => 32767,
    1450 => 32767,
    1451 => 32767,
    1452 => 32767,
    1453 => 32767,
    1454 => 32767,
    1455 => 32767,
    1456 => 32767,
    1457 => 32767,
    1458 => 32767,
    1459 => 32767,
    1460 => 32767,
    1461 => 32767,
    1462 => 32767,
    1463 => 32767,
    1464 => 32767,
    1465 => 32767,
    1466 => 32767,
    1467 => 32767,
    1468 => 32767,
    1469 => 32767,
    1470 => 32767,
    1471 => 32767,
    1472 => 32767,
    1473 => 32767,
    1474 => 32767,
    1475 => 32767,
    1476 => 32767,
    1477 => 32767,
    1478 => 32767,
    1479 => 32767,
    1480 => 32767,
    1481 => 32767,
    1482 => 32767,
    1483 => 32767,
    1484 => 32767,
    1485 => 32767,
    1486 => 32767,
    1487 => 32767,
    1488 => 32767,
    1489 => 32767,
    1490 => 32767,
    1491 => 32767,
    1492 => 32767,
    1493 => 32767,
    1494 => 32767,
    1495 => 32767,
    1496 => 32767,
    1497 => 32767,
    1498 => 32767,
    1499 => 32767,
    1500 => 32767,
    1501 => 32767,
    1502 => 32767,
    1503 => 32767,
    1504 => 32767,
    1505 => 32767,
    1506 => 32767,
    1507 => 32767,
    1508 => 32767,
    1509 => 32767,
    1510 => 32767,
    1511 => 32767,
    1512 => 32767,
    1513 => 32767,
    1514 => 32767,
    1515 => 32767,
    1516 => 32767,
    1517 => 32767,
    1518 => 32767,
    1519 => 32767,
    1520 => 32767,
    1521 => 32767,
    1522 => 32767,
    1523 => 32767,
    1524 => 32767,
    1525 => 32767,
    1526 => 32767,
    1527 => 32767,
    1528 => 32767,
    1529 => 32767,
    1530 => 32767,
    1531 => 32767,
    1532 => 32767,
    1533 => 32767,
    1534 => 32767,
    1535 => 32767,
    1536 => 32767,
    1537 => 32767,
    1538 => 32767,
    1539 => 32767,
    1540 => 32767,
    1541 => 32767,
    1542 => 32767,
    1543 => 32767,
    1544 => 32767,
    1545 => 32767,
    1546 => 32767,
    1547 => 32767,
    1548 => 32767,
    1549 => 32767,
    1550 => 32767,
    1551 => 32767,
    1552 => 32767,
    1553 => 32767,
    1554 => 32767,
    1555 => 32767,
    1556 => 32767,
    1557 => 32767,
    1558 => 32767,
    1559 => 32767,
    1560 => 32767,
    1561 => 32767,
    1562 => 32767,
    1563 => 32767,
    1564 => 32767,
    1565 => 32767,
    1566 => 32767,
    1567 => 32767,
    1568 => 32767,
    1569 => 32767,
    1570 => 32767,
    1571 => 32767,
    1572 => 32767,
    1573 => 32767,
    1574 => 32767,
    1575 => 32767,
    1576 => 32767,
    1577 => 32767,
    1578 => 32767,
    1579 => 32767,
    1580 => 32767,
    1581 => 32767,
    1582 => 32767,
    1583 => 32767,
    1584 => 32767,
    1585 => 32767,
    1586 => 32767,
    1587 => 32767,
    1588 => 32767,
    1589 => 32767,
    1590 => 32767,
    1591 => 32767,
    1592 => 32767,
    1593 => 32767,
    1594 => 32767,
    1595 => 32767,
    1596 => 32767,
    1597 => 32767,
    1598 => 32767,
    1599 => 32767,
    1600 => 32767,
    1601 => 32767,
    1602 => 32767,
    1603 => 32767,
    1604 => 32767,
    1605 => 32767,
    1606 => 32767,
    1607 => 32767,
    1608 => 32767,
    1609 => 32767,
    1610 => 32767,
    1611 => 32767,
    1612 => 32767,
    1613 => 32767,
    1614 => 32767,
    1615 => 32767,
    1616 => 32767,
    1617 => 32767,
    1618 => 32767,
    1619 => 32767,
    1620 => 32767,
    1621 => 32767,
    1622 => 32767,
    1623 => 32767,
    1624 => 32767,
    1625 => 32767,
    1626 => 32767,
    1627 => 32767,
    1628 => 32767,
    1629 => 32767,
    1630 => 32767,
    1631 => 32767,
    1632 => 32767,
    1633 => 32767,
    1634 => 32767,
    1635 => 32767,
    1636 => 32767,
    1637 => 32767,
    1638 => 32767,
    1639 => 32767,
    1640 => 32767,
    1641 => 32767,
    1642 => 32767,
    1643 => 32767,
    1644 => 32767,
    1645 => 32767,
    1646 => 32767,
    1647 => 32767,
    1648 => 32767,
    1649 => 32767,
    1650 => 32767,
    1651 => 32767,
    1652 => 32767,
    1653 => 32767,
    1654 => 32767,
    1655 => 32767,
    1656 => 32767,
    1657 => 32767,
    1658 => 32767,
    1659 => 32767,
    1660 => 32767,
    1661 => 32767,
    1662 => 32767,
    1663 => 32767,
    1664 => 32767,
    1665 => 32767,
    1666 => 32767,
    1667 => 32767,
    1668 => 32767,
    1669 => 32767,
    1670 => 32767,
    1671 => 32767,
    1672 => 32767,
    1673 => 32767,
    1674 => 32767,
    1675 => 32767,
    1676 => 32767,
    1677 => 32767,
    1678 => 32767,
    1679 => 32767,
    1680 => 32767,
    1681 => 32767,
    1682 => 32767,
    1683 => 32767,
    1684 => 32767,
    1685 => 32767,
    1686 => 32767,
    1687 => 32767,
    1688 => 32767,
    1689 => 32767,
    1690 => 32767,
    1691 => 32767,
    1692 => 32767,
    1693 => 32767,
    1694 => 32767,
    1695 => 32767,
    1696 => 32767,
    1697 => 32767,
    1698 => 32767,
    1699 => 32767,
    1700 => 32767,
    1701 => 32767,
    1702 => 32767,
    1703 => 32767,
    1704 => 32767,
    1705 => 32767,
    1706 => 32767,
    1707 => 32767,
    1708 => 32767,
    1709 => 32767,
    1710 => 32767,
    1711 => 32767,
    1712 => 32767,
    1713 => 32767,
    1714 => 32767,
    1715 => 32767,
    1716 => 32767,
    1717 => 32767,
    1718 => 32767,
    1719 => 32767,
    1720 => 32767,
    1721 => 32767,
    1722 => 32767,
    1723 => 32767,
    1724 => 32767,
    1725 => 32767,
    1726 => 32767,
    1727 => 32767,
    1728 => 32767,
    1729 => 32767,
    1730 => 32767,
    1731 => 32767,
    1732 => 32767,
    1733 => 32767,
    1734 => 32767,
    1735 => 32767,
    1736 => 32767,
    1737 => 32767,
    1738 => 32767,
    1739 => 32767,
    1740 => 32767,
    1741 => 32767,
    1742 => 32767,
    1743 => 32767,
    1744 => 32767,
    1745 => 32767,
    1746 => 32767,
    1747 => 32767,
    1748 => 32767,
    1749 => 32767,
    1750 => 32767,
    1751 => 32767,
    1752 => 32767,
    1753 => 32767,
    1754 => 32767,
    1755 => 32767,
    1756 => 32767,
    1757 => 32767,
    1758 => 32767,
    1759 => 32767,
    1760 => 32767,
    1761 => 32767,
    1762 => 32767,
    1763 => 32767,
    1764 => 32767,
    1765 => 32767,
    1766 => 32767,
    1767 => 32767,
    1768 => 32767,
    1769 => 32767,
    1770 => 32767,
    1771 => 32767,
    1772 => 32767,
    1773 => 32767,
    1774 => 32767,
    1775 => 32767,
    1776 => 32767,
    1777 => 32767,
    1778 => 32767,
    1779 => 32767,
    1780 => 32767,
    1781 => 32767,
    1782 => 32767,
    1783 => 32767,
    1784 => 32767,
    1785 => 32767,
    1786 => 32767,
    1787 => 32767,
    1788 => 32767,
    1789 => 32767,
    1790 => 32767,
    1791 => 32767,
    1792 => 32767,
    1793 => 32767,
    1794 => 32767,
    1795 => 32767,
    1796 => 32767,
    1797 => 32767,
    1798 => 32767,
    1799 => 32767,
    1800 => 32767,
    1801 => 32767,
    1802 => 32767,
    1803 => 32767,
    1804 => 32767,
    1805 => 32767,
    1806 => 32767,
    1807 => 32767,
    1808 => 32767,
    1809 => 32767,
    1810 => 32767,
    1811 => 32767,
    1812 => 32767,
    1813 => 32767,
    1814 => 32767,
    1815 => 32767,
    1816 => 32767,
    1817 => 32767,
    1818 => 32767,
    1819 => 32767,
    1820 => 32767,
    1821 => 32767,
    1822 => 32767,
    1823 => 32767,
    1824 => 32767,
    1825 => 32767,
    1826 => 32767,
    1827 => 32767,
    1828 => 32767,
    1829 => 32767,
    1830 => 32767,
    1831 => 32767,
    1832 => 32767,
    1833 => 32767,
    1834 => 32767,
    1835 => 32767,
    1836 => 32767,
    1837 => 32767,
    1838 => 32767,
    1839 => 32767,
    1840 => 32767,
    1841 => 32767,
    1842 => 32767,
    1843 => 32767,
    1844 => 32767,
    1845 => 32767,
    1846 => 32767,
    1847 => 32767,
    1848 => 32767,
    1849 => 32767,
    1850 => 32767,
    1851 => 32767,
    1852 => 32767,
    1853 => 32767,
    1854 => 32767,
    1855 => 32767,
    1856 => 32767,
    1857 => 32767,
    1858 => 32767,
    1859 => 32767,
    1860 => 32767,
    1861 => 32767,
    1862 => 32767,
    1863 => 32767,
    1864 => 32767,
    1865 => 32767,
    1866 => 32767,
    1867 => 32767,
    1868 => 32767,
    1869 => 32767,
    1870 => 32767,
    1871 => 32767,
    1872 => 32767,
    1873 => 32767,
    1874 => 32767,
    1875 => 32767,
    1876 => 32767,
    1877 => 32767,
    1878 => 32767,
    1879 => 32767,
    1880 => 32767,
    1881 => 32767,
    1882 => 32767,
    1883 => 32767,
    1884 => 32767,
    1885 => 32767,
    1886 => 32767,
    1887 => 32767,
    1888 => 32767,
    1889 => 32767,
    1890 => 32767,
    1891 => 32767,
    1892 => 32767,
    1893 => 32767,
    1894 => 32767,
    1895 => 32767,
    1896 => 32767,
    1897 => 32767,
    1898 => 32767,
    1899 => 32767,
    1900 => 32767,
    1901 => 32767,
    1902 => 32767,
    1903 => 32767,
    1904 => 32767,
    1905 => 32767,
    1906 => 32767,
    1907 => 32767,
    1908 => 32767,
    1909 => 32767,
    1910 => 32767,
    1911 => 32767,
    1912 => 32767,
    1913 => 32767,
    1914 => 32767,
    1915 => 32767,
    1916 => 32767,
    1917 => 32767,
    1918 => 32767,
    1919 => 32767,
    1920 => 32767,
    1921 => 32767,
    1922 => 32767,
    1923 => 32767,
    1924 => 32767,
    1925 => 32767,
    1926 => 32767,
    1927 => 32767,
    1928 => 32767,
    1929 => 32767,
    1930 => 32767,
    1931 => 32767,
    1932 => 32767,
    1933 => 32767,
    1934 => 32767,
    1935 => 32767,
    1936 => 32767,
    1937 => 32767,
    1938 => 32767,
    1939 => 32767,
    1940 => 32767,
    1941 => 32767,
    1942 => 32767,
    1943 => 32767,
    1944 => 32767,
    1945 => 32767,
    1946 => 32767,
    1947 => 32767,
    1948 => 32767,
    1949 => 32767,
    1950 => 32767,
    1951 => 32767,
    1952 => 32767,
    1953 => 32767,
    1954 => 32767,
    1955 => 32767,
    1956 => 32767,
    1957 => 32767,
    1958 => 32767,
    1959 => 32767,
    1960 => 32767,
    1961 => 32767,
    1962 => 32767,
    1963 => 32767,
    1964 => 32767,
    1965 => 32767,
    1966 => 32767,
    1967 => 32767,
    1968 => 32767,
    1969 => 32767,
    1970 => 32767,
    1971 => 32767,
    1972 => 32767,
    1973 => 32767,
    1974 => 32767,
    1975 => 32767,
    1976 => 32767,
    1977 => 32767,
    1978 => 32767,
    1979 => 32767,
    1980 => 32767,
    1981 => 32767,
    1982 => 32767,
    1983 => 32767,
    1984 => 32767,
    1985 => 32767,
    1986 => 32767,
    1987 => 32767,
    1988 => 32767,
    1989 => 32767,
    1990 => 32767,
    1991 => 32767,
    1992 => 32767,
    1993 => 32767,
    1994 => 32767,
    1995 => 32767,
    1996 => 32767,
    1997 => 32767,
    1998 => 32767,
    1999 => 32767,
    2000 => 32767,
    2001 => 32767,
    2002 => 32767,
    2003 => 32767,
    2004 => 32767,
    2005 => 32767,
    2006 => 32767,
    2007 => 32767,
    2008 => 32767,
    2009 => 32767,
    2010 => 32767,
    2011 => 32767,
    2012 => 32767,
    2013 => 32767,
    2014 => 32767,
    2015 => 32767,
    2016 => 32767,
    2017 => 32767,
    2018 => 32767,
    2019 => 32767,
    2020 => 32767,
    2021 => 32767,
    2022 => 32767,
    2023 => 32767,
    2024 => 32767,
    2025 => 32767,
    2026 => 32767,
    2027 => 32767,
    2028 => 32767,
    2029 => 32767,
    2030 => 32767,
    2031 => 32767,
    2032 => 32767,
    2033 => 32767,
    2034 => 32767,
    2035 => 32767,
    2036 => 32767,
    2037 => 32767,
    2038 => 32767,
    2039 => 32767,
    2040 => 32767,
    2041 => 32767,
    2042 => 32767,
    2043 => 32767,
    2044 => 32767,
    2045 => 32767,
    2046 => 32767,
    2047 => 32767
);

begin
  dds_out <= std_logic_vector(TO_SIGNED(LUT(TO_INTEGER(unsigned(address))),16));
end rtl;
