library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sigmoid_lut_2048 is
  port (
    address : in  std_logic_vector(11 downto 0);
    dds_out : out std_logic_vector(15 downto 0) 
  );
end sigmoid_lut_2048;


-- Output between [-11; +11], rapresented with fixed point
-- Need for 1 bit for integer, last 15 bit for float rapresentation
-- Reach the LSB method
-- 
-- LSB(in) = (11)/(2^11 - 1) = 0.00537371763556424035173424523693
-- LSB(out) = (1)/(2^15 - 1) = 3.0518509475997192297128208258309e-5
-- inputs -> [-11, +11] 
-- outputs -> [0, 1]
-- Q(f(x)) = round(f(x)/LSB(out))*LSB(out)
-- 
--
-- What to store in the lut? round(f(x)/LSB(out)) for x in [0; 2047]*LSB(in)

architecture rtl of sigmoid_lut_2048 is
type LUT_t is array (natural range 0 to 2047) of integer;
constant LUT: LUT_t := (
    0 => 16384,
    1 => 16428,
    2 => 16472,
    3 => 16516,
    4 => 16560,
    5 => 16604,
    6 => 16648,
    7 => 16692,
    8 => 16736,
    9 => 16780,
    10 => 16824,
    11 => 16868,
    12 => 16912,
    13 => 16956,
    14 => 16999,
    15 => 17043,
    16 => 17087,
    17 => 17131,
    18 => 17175,
    19 => 17219,
    20 => 17263,
    21 => 17307,
    22 => 17351,
    23 => 17395,
    24 => 17439,
    25 => 17482,
    26 => 17526,
    27 => 17570,
    28 => 17614,
    29 => 17658,
    30 => 17701,
    31 => 17745,
    32 => 17789,
    33 => 17832,
    34 => 17876,
    35 => 17920,
    36 => 17963,
    37 => 18007,
    38 => 18050,
    39 => 18094,
    40 => 18138,
    41 => 18181,
    42 => 18225,
    43 => 18268,
    44 => 18311,
    45 => 18355,
    46 => 18398,
    47 => 18442,
    48 => 18485,
    49 => 18528,
    50 => 18571,
    51 => 18615,
    52 => 18658,
    53 => 18701,
    54 => 18744,
    55 => 18787,
    56 => 18830,
    57 => 18873,
    58 => 18916,
    59 => 18959,
    60 => 19002,
    61 => 19045,
    62 => 19088,
    63 => 19131,
    64 => 19173,
    65 => 19216,
    66 => 19259,
    67 => 19301,
    68 => 19344,
    69 => 19387,
    70 => 19429,
    71 => 19472,
    72 => 19514,
    73 => 19556,
    74 => 19599,
    75 => 19641,
    76 => 19683,
    77 => 19726,
    78 => 19768,
    79 => 19810,
    80 => 19852,
    81 => 19894,
    82 => 19936,
    83 => 19978,
    84 => 20020,
    85 => 20061,
    86 => 20103,
    87 => 20145,
    88 => 20187,
    89 => 20228,
    90 => 20270,
    91 => 20311,
    92 => 20353,
    93 => 20394,
    94 => 20436,
    95 => 20477,
    96 => 20518,
    97 => 20559,
    98 => 20600,
    99 => 20642,
    100 => 20683,
    101 => 20724,
    102 => 20764,
    103 => 20805,
    104 => 20846,
    105 => 20887,
    106 => 20927,
    107 => 20968,
    108 => 21009,
    109 => 21049,
    110 => 21089,
    111 => 21130,
    112 => 21170,
    113 => 21210,
    114 => 21251,
    115 => 21291,
    116 => 21331,
    117 => 21371,
    118 => 21411,
    119 => 21450,
    120 => 21490,
    121 => 21530,
    122 => 21570,
    123 => 21609,
    124 => 21649,
    125 => 21688,
    126 => 21727,
    127 => 21767,
    128 => 21806,
    129 => 21845,
    130 => 21884,
    131 => 21923,
    132 => 21962,
    133 => 22001,
    134 => 22040,
    135 => 22079,
    136 => 22117,
    137 => 22156,
    138 => 22194,
    139 => 22233,
    140 => 22271,
    141 => 22310,
    142 => 22348,
    143 => 22386,
    144 => 22424,
    145 => 22462,
    146 => 22500,
    147 => 22538,
    148 => 22575,
    149 => 22613,
    150 => 22651,
    151 => 22688,
    152 => 22726,
    153 => 22763,
    154 => 22800,
    155 => 22838,
    156 => 22875,
    157 => 22912,
    158 => 22949,
    159 => 22986,
    160 => 23023,
    161 => 23059,
    162 => 23096,
    163 => 23133,
    164 => 23169,
    165 => 23206,
    166 => 23242,
    167 => 23278,
    168 => 23314,
    169 => 23351,
    170 => 23387,
    171 => 23422,
    172 => 23458,
    173 => 23494,
    174 => 23530,
    175 => 23565,
    176 => 23601,
    177 => 23636,
    178 => 23672,
    179 => 23707,
    180 => 23742,
    181 => 23777,
    182 => 23812,
    183 => 23847,
    184 => 23882,
    185 => 23917,
    186 => 23951,
    187 => 23986,
    188 => 24021,
    189 => 24055,
    190 => 24089,
    191 => 24124,
    192 => 24158,
    193 => 24192,
    194 => 24226,
    195 => 24260,
    196 => 24293,
    197 => 24327,
    198 => 24361,
    199 => 24394,
    200 => 24428,
    201 => 24461,
    202 => 24494,
    203 => 24528,
    204 => 24561,
    205 => 24594,
    206 => 24627,
    207 => 24659,
    208 => 24692,
    209 => 24725,
    210 => 24757,
    211 => 24790,
    212 => 24822,
    213 => 24855,
    214 => 24887,
    215 => 24919,
    216 => 24951,
    217 => 24983,
    218 => 25015,
    219 => 25046,
    220 => 25078,
    221 => 25110,
    222 => 25141,
    223 => 25173,
    224 => 25204,
    225 => 25235,
    226 => 25266,
    227 => 25297,
    228 => 25328,
    229 => 25359,
    230 => 25390,
    231 => 25420,
    232 => 25451,
    233 => 25482,
    234 => 25512,
    235 => 25542,
    236 => 25572,
    237 => 25603,
    238 => 25633,
    239 => 25663,
    240 => 25692,
    241 => 25722,
    242 => 25752,
    243 => 25781,
    244 => 25811,
    245 => 25840,
    246 => 25870,
    247 => 25899,
    248 => 25928,
    249 => 25957,
    250 => 25986,
    251 => 26015,
    252 => 26044,
    253 => 26072,
    254 => 26101,
    255 => 26129,
    256 => 26158,
    257 => 26186,
    258 => 26214,
    259 => 26242,
    260 => 26270,
    261 => 26298,
    262 => 26326,
    263 => 26354,
    264 => 26382,
    265 => 26409,
    266 => 26437,
    267 => 26464,
    268 => 26491,
    269 => 26519,
    270 => 26546,
    271 => 26573,
    272 => 26600,
    273 => 26627,
    274 => 26653,
    275 => 26680,
    276 => 26707,
    277 => 26733,
    278 => 26760,
    279 => 26786,
    280 => 26812,
    281 => 26838,
    282 => 26864,
    283 => 26890,
    284 => 26916,
    285 => 26942,
    286 => 26968,
    287 => 26993,
    288 => 27019,
    289 => 27044,
    290 => 27069,
    291 => 27095,
    292 => 27120,
    293 => 27145,
    294 => 27170,
    295 => 27195,
    296 => 27220,
    297 => 27244,
    298 => 27269,
    299 => 27294,
    300 => 27318,
    301 => 27342,
    302 => 27367,
    303 => 27391,
    304 => 27415,
    305 => 27439,
    306 => 27463,
    307 => 27487,
    308 => 27511,
    309 => 27534,
    310 => 27558,
    311 => 27581,
    312 => 27605,
    313 => 27628,
    314 => 27651,
    315 => 27674,
    316 => 27697,
    317 => 27720,
    318 => 27743,
    319 => 27766,
    320 => 27789,
    321 => 27812,
    322 => 27834,
    323 => 27857,
    324 => 27879,
    325 => 27901,
    326 => 27924,
    327 => 27946,
    328 => 27968,
    329 => 27990,
    330 => 28012,
    331 => 28033,
    332 => 28055,
    333 => 28077,
    334 => 28098,
    335 => 28120,
    336 => 28141,
    337 => 28162,
    338 => 28184,
    339 => 28205,
    340 => 28226,
    341 => 28247,
    342 => 28268,
    343 => 28289,
    344 => 28309,
    345 => 28330,
    346 => 28351,
    347 => 28371,
    348 => 28391,
    349 => 28412,
    350 => 28432,
    351 => 28452,
    352 => 28472,
    353 => 28492,
    354 => 28512,
    355 => 28532,
    356 => 28552,
    357 => 28572,
    358 => 28591,
    359 => 28611,
    360 => 28630,
    361 => 28650,
    362 => 28669,
    363 => 28688,
    364 => 28707,
    365 => 28726,
    366 => 28745,
    367 => 28764,
    368 => 28783,
    369 => 28802,
    370 => 28821,
    371 => 28839,
    372 => 28858,
    373 => 28876,
    374 => 28895,
    375 => 28913,
    376 => 28931,
    377 => 28949,
    378 => 28967,
    379 => 28985,
    380 => 29003,
    381 => 29021,
    382 => 29039,
    383 => 29057,
    384 => 29074,
    385 => 29092,
    386 => 29109,
    387 => 29127,
    388 => 29144,
    389 => 29161,
    390 => 29179,
    391 => 29196,
    392 => 29213,
    393 => 29230,
    394 => 29247,
    395 => 29264,
    396 => 29280,
    397 => 29297,
    398 => 29314,
    399 => 29330,
    400 => 29347,
    401 => 29363,
    402 => 29380,
    403 => 29396,
    404 => 29412,
    405 => 29428,
    406 => 29444,
    407 => 29460,
    408 => 29476,
    409 => 29492,
    410 => 29508,
    411 => 29524,
    412 => 29539,
    413 => 29555,
    414 => 29570,
    415 => 29586,
    416 => 29601,
    417 => 29617,
    418 => 29632,
    419 => 29647,
    420 => 29662,
    421 => 29677,
    422 => 29692,
    423 => 29707,
    424 => 29722,
    425 => 29737,
    426 => 29752,
    427 => 29766,
    428 => 29781,
    429 => 29796,
    430 => 29810,
    431 => 29825,
    432 => 29839,
    433 => 29853,
    434 => 29867,
    435 => 29882,
    436 => 29896,
    437 => 29910,
    438 => 29924,
    439 => 29938,
    440 => 29951,
    441 => 29965,
    442 => 29979,
    443 => 29993,
    444 => 30006,
    445 => 30020,
    446 => 30033,
    447 => 30047,
    448 => 30060,
    449 => 30073,
    450 => 30087,
    451 => 30100,
    452 => 30113,
    453 => 30126,
    454 => 30139,
    455 => 30152,
    456 => 30165,
    457 => 30178,
    458 => 30191,
    459 => 30203,
    460 => 30216,
    461 => 30229,
    462 => 30241,
    463 => 30254,
    464 => 30266,
    465 => 30279,
    466 => 30291,
    467 => 30303,
    468 => 30315,
    469 => 30328,
    470 => 30340,
    471 => 30352,
    472 => 30364,
    473 => 30376,
    474 => 30388,
    475 => 30399,
    476 => 30411,
    477 => 30423,
    478 => 30435,
    479 => 30446,
    480 => 30458,
    481 => 30469,
    482 => 30481,
    483 => 30492,
    484 => 30503,
    485 => 30515,
    486 => 30526,
    487 => 30537,
    488 => 30548,
    489 => 30559,
    490 => 30570,
    491 => 30581,
    492 => 30592,
    493 => 30603,
    494 => 30614,
    495 => 30625,
    496 => 30636,
    497 => 30646,
    498 => 30657,
    499 => 30667,
    500 => 30678,
    501 => 30688,
    502 => 30699,
    503 => 30709,
    504 => 30720,
    505 => 30730,
    506 => 30740,
    507 => 30750,
    508 => 30761,
    509 => 30771,
    510 => 30781,
    511 => 30791,
    512 => 30801,
    513 => 30811,
    514 => 30820,
    515 => 30830,
    516 => 30840,
    517 => 30850,
    518 => 30859,
    519 => 30869,
    520 => 30879,
    521 => 30888,
    522 => 30898,
    523 => 30907,
    524 => 30916,
    525 => 30926,
    526 => 30935,
    527 => 30944,
    528 => 30954,
    529 => 30963,
    530 => 30972,
    531 => 30981,
    532 => 30990,
    533 => 30999,
    534 => 31008,
    535 => 31017,
    536 => 31026,
    537 => 31035,
    538 => 31044,
    539 => 31052,
    540 => 31061,
    541 => 31070,
    542 => 31078,
    543 => 31087,
    544 => 31095,
    545 => 31104,
    546 => 31112,
    547 => 31121,
    548 => 31129,
    549 => 31138,
    550 => 31146,
    551 => 31154,
    552 => 31162,
    553 => 31171,
    554 => 31179,
    555 => 31187,
    556 => 31195,
    557 => 31203,
    558 => 31211,
    559 => 31219,
    560 => 31227,
    561 => 31235,
    562 => 31242,
    563 => 31250,
    564 => 31258,
    565 => 31266,
    566 => 31273,
    567 => 31281,
    568 => 31289,
    569 => 31296,
    570 => 31304,
    571 => 31311,
    572 => 31319,
    573 => 31326,
    574 => 31333,
    575 => 31341,
    576 => 31348,
    577 => 31355,
    578 => 31363,
    579 => 31370,
    580 => 31377,
    581 => 31384,
    582 => 31391,
    583 => 31398,
    584 => 31405,
    585 => 31412,
    586 => 31419,
    587 => 31426,
    588 => 31433,
    589 => 31440,
    590 => 31447,
    591 => 31454,
    592 => 31460,
    593 => 31467,
    594 => 31474,
    595 => 31480,
    596 => 31487,
    597 => 31494,
    598 => 31500,
    599 => 31507,
    600 => 31513,
    601 => 31520,
    602 => 31526,
    603 => 31532,
    604 => 31539,
    605 => 31545,
    606 => 31552,
    607 => 31558,
    608 => 31564,
    609 => 31570,
    610 => 31576,
    611 => 31583,
    612 => 31589,
    613 => 31595,
    614 => 31601,
    615 => 31607,
    616 => 31613,
    617 => 31619,
    618 => 31625,
    619 => 31631,
    620 => 31637,
    621 => 31642,
    622 => 31648,
    623 => 31654,
    624 => 31660,
    625 => 31666,
    626 => 31671,
    627 => 31677,
    628 => 31683,
    629 => 31688,
    630 => 31694,
    631 => 31699,
    632 => 31705,
    633 => 31710,
    634 => 31716,
    635 => 31721,
    636 => 31727,
    637 => 31732,
    638 => 31738,
    639 => 31743,
    640 => 31748,
    641 => 31753,
    642 => 31759,
    643 => 31764,
    644 => 31769,
    645 => 31774,
    646 => 31780,
    647 => 31785,
    648 => 31790,
    649 => 31795,
    650 => 31800,
    651 => 31805,
    652 => 31810,
    653 => 31815,
    654 => 31820,
    655 => 31825,
    656 => 31830,
    657 => 31835,
    658 => 31839,
    659 => 31844,
    660 => 31849,
    661 => 31854,
    662 => 31859,
    663 => 31863,
    664 => 31868,
    665 => 31873,
    666 => 31877,
    667 => 31882,
    668 => 31887,
    669 => 31891,
    670 => 31896,
    671 => 31900,
    672 => 31905,
    673 => 31909,
    674 => 31914,
    675 => 31918,
    676 => 31923,
    677 => 31927,
    678 => 31932,
    679 => 31936,
    680 => 31940,
    681 => 31945,
    682 => 31949,
    683 => 31953,
    684 => 31957,
    685 => 31962,
    686 => 31966,
    687 => 31970,
    688 => 31974,
    689 => 31978,
    690 => 31982,
    691 => 31987,
    692 => 31991,
    693 => 31995,
    694 => 31999,
    695 => 32003,
    696 => 32007,
    697 => 32011,
    698 => 32015,
    699 => 32019,
    700 => 32023,
    701 => 32026,
    702 => 32030,
    703 => 32034,
    704 => 32038,
    705 => 32042,
    706 => 32046,
    707 => 32049,
    708 => 32053,
    709 => 32057,
    710 => 32061,
    711 => 32064,
    712 => 32068,
    713 => 32072,
    714 => 32075,
    715 => 32079,
    716 => 32083,
    717 => 32086,
    718 => 32090,
    719 => 32093,
    720 => 32097,
    721 => 32100,
    722 => 32104,
    723 => 32107,
    724 => 32111,
    725 => 32114,
    726 => 32118,
    727 => 32121,
    728 => 32125,
    729 => 32128,
    730 => 32131,
    731 => 32135,
    732 => 32138,
    733 => 32141,
    734 => 32145,
    735 => 32148,
    736 => 32151,
    737 => 32154,
    738 => 32158,
    739 => 32161,
    740 => 32164,
    741 => 32167,
    742 => 32170,
    743 => 32173,
    744 => 32177,
    745 => 32180,
    746 => 32183,
    747 => 32186,
    748 => 32189,
    749 => 32192,
    750 => 32195,
    751 => 32198,
    752 => 32201,
    753 => 32204,
    754 => 32207,
    755 => 32210,
    756 => 32213,
    757 => 32216,
    758 => 32219,
    759 => 32221,
    760 => 32224,
    761 => 32227,
    762 => 32230,
    763 => 32233,
    764 => 32236,
    765 => 32239,
    766 => 32241,
    767 => 32244,
    768 => 32247,
    769 => 32250,
    770 => 32252,
    771 => 32255,
    772 => 32258,
    773 => 32260,
    774 => 32263,
    775 => 32266,
    776 => 32268,
    777 => 32271,
    778 => 32274,
    779 => 32276,
    780 => 32279,
    781 => 32281,
    782 => 32284,
    783 => 32287,
    784 => 32289,
    785 => 32292,
    786 => 32294,
    787 => 32297,
    788 => 32299,
    789 => 32302,
    790 => 32304,
    791 => 32306,
    792 => 32309,
    793 => 32311,
    794 => 32314,
    795 => 32316,
    796 => 32318,
    797 => 32321,
    798 => 32323,
    799 => 32326,
    800 => 32328,
    801 => 32330,
    802 => 32333,
    803 => 32335,
    804 => 32337,
    805 => 32339,
    806 => 32342,
    807 => 32344,
    808 => 32346,
    809 => 32348,
    810 => 32351,
    811 => 32353,
    812 => 32355,
    813 => 32357,
    814 => 32359,
    815 => 32361,
    816 => 32364,
    817 => 32366,
    818 => 32368,
    819 => 32370,
    820 => 32372,
    821 => 32374,
    822 => 32376,
    823 => 32378,
    824 => 32380,
    825 => 32382,
    826 => 32384,
    827 => 32387,
    828 => 32389,
    829 => 32391,
    830 => 32393,
    831 => 32395,
    832 => 32396,
    833 => 32398,
    834 => 32400,
    835 => 32402,
    836 => 32404,
    837 => 32406,
    838 => 32408,
    839 => 32410,
    840 => 32412,
    841 => 32414,
    842 => 32416,
    843 => 32418,
    844 => 32419,
    845 => 32421,
    846 => 32423,
    847 => 32425,
    848 => 32427,
    849 => 32429,
    850 => 32430,
    851 => 32432,
    852 => 32434,
    853 => 32436,
    854 => 32437,
    855 => 32439,
    856 => 32441,
    857 => 32443,
    858 => 32444,
    859 => 32446,
    860 => 32448,
    861 => 32449,
    862 => 32451,
    863 => 32453,
    864 => 32454,
    865 => 32456,
    866 => 32458,
    867 => 32459,
    868 => 32461,
    869 => 32463,
    870 => 32464,
    871 => 32466,
    872 => 32468,
    873 => 32469,
    874 => 32471,
    875 => 32472,
    876 => 32474,
    877 => 32475,
    878 => 32477,
    879 => 32478,
    880 => 32480,
    881 => 32482,
    882 => 32483,
    883 => 32485,
    884 => 32486,
    885 => 32488,
    886 => 32489,
    887 => 32490,
    888 => 32492,
    889 => 32493,
    890 => 32495,
    891 => 32496,
    892 => 32498,
    893 => 32499,
    894 => 32501,
    895 => 32502,
    896 => 32503,
    897 => 32505,
    898 => 32506,
    899 => 32508,
    900 => 32509,
    901 => 32510,
    902 => 32512,
    903 => 32513,
    904 => 32514,
    905 => 32516,
    906 => 32517,
    907 => 32518,
    908 => 32520,
    909 => 32521,
    910 => 32522,
    911 => 32524,
    912 => 32525,
    913 => 32526,
    914 => 32528,
    915 => 32529,
    916 => 32530,
    917 => 32531,
    918 => 32533,
    919 => 32534,
    920 => 32535,
    921 => 32536,
    922 => 32538,
    923 => 32539,
    924 => 32540,
    925 => 32541,
    926 => 32542,
    927 => 32544,
    928 => 32545,
    929 => 32546,
    930 => 32547,
    931 => 32548,
    932 => 32549,
    933 => 32551,
    934 => 32552,
    935 => 32553,
    936 => 32554,
    937 => 32555,
    938 => 32556,
    939 => 32557,
    940 => 32559,
    941 => 32560,
    942 => 32561,
    943 => 32562,
    944 => 32563,
    945 => 32564,
    946 => 32565,
    947 => 32566,
    948 => 32567,
    949 => 32568,
    950 => 32569,
    951 => 32570,
    952 => 32572,
    953 => 32573,
    954 => 32574,
    955 => 32575,
    956 => 32576,
    957 => 32577,
    958 => 32578,
    959 => 32579,
    960 => 32580,
    961 => 32581,
    962 => 32582,
    963 => 32583,
    964 => 32584,
    965 => 32585,
    966 => 32586,
    967 => 32587,
    968 => 32588,
    969 => 32589,
    970 => 32589,
    971 => 32590,
    972 => 32591,
    973 => 32592,
    974 => 32593,
    975 => 32594,
    976 => 32595,
    977 => 32596,
    978 => 32597,
    979 => 32598,
    980 => 32599,
    981 => 32600,
    982 => 32600,
    983 => 32601,
    984 => 32602,
    985 => 32603,
    986 => 32604,
    987 => 32605,
    988 => 32606,
    989 => 32607,
    990 => 32607,
    991 => 32608,
    992 => 32609,
    993 => 32610,
    994 => 32611,
    995 => 32612,
    996 => 32612,
    997 => 32613,
    998 => 32614,
    999 => 32615,
    1000 => 32616,
    1001 => 32617,
    1002 => 32617,
    1003 => 32618,
    1004 => 32619,
    1005 => 32620,
    1006 => 32621,
    1007 => 32621,
    1008 => 32622,
    1009 => 32623,
    1010 => 32624,
    1011 => 32624,
    1012 => 32625,
    1013 => 32626,
    1014 => 32627,
    1015 => 32627,
    1016 => 32628,
    1017 => 32629,
    1018 => 32630,
    1019 => 32630,
    1020 => 32631,
    1021 => 32632,
    1022 => 32633,
    1023 => 32633,
    1024 => 32634,
    1025 => 32635,
    1026 => 32635,
    1027 => 32636,
    1028 => 32637,
    1029 => 32638,
    1030 => 32638,
    1031 => 32639,
    1032 => 32640,
    1033 => 32640,
    1034 => 32641,
    1035 => 32642,
    1036 => 32642,
    1037 => 32643,
    1038 => 32644,
    1039 => 32644,
    1040 => 32645,
    1041 => 32646,
    1042 => 32646,
    1043 => 32647,
    1044 => 32647,
    1045 => 32648,
    1046 => 32649,
    1047 => 32649,
    1048 => 32650,
    1049 => 32651,
    1050 => 32651,
    1051 => 32652,
    1052 => 32653,
    1053 => 32653,
    1054 => 32654,
    1055 => 32654,
    1056 => 32655,
    1057 => 32656,
    1058 => 32656,
    1059 => 32657,
    1060 => 32657,
    1061 => 32658,
    1062 => 32658,
    1063 => 32659,
    1064 => 32660,
    1065 => 32660,
    1066 => 32661,
    1067 => 32661,
    1068 => 32662,
    1069 => 32662,
    1070 => 32663,
    1071 => 32664,
    1072 => 32664,
    1073 => 32665,
    1074 => 32665,
    1075 => 32666,
    1076 => 32666,
    1077 => 32667,
    1078 => 32667,
    1079 => 32668,
    1080 => 32668,
    1081 => 32669,
    1082 => 32670,
    1083 => 32670,
    1084 => 32671,
    1085 => 32671,
    1086 => 32672,
    1087 => 32672,
    1088 => 32673,
    1089 => 32673,
    1090 => 32674,
    1091 => 32674,
    1092 => 32675,
    1093 => 32675,
    1094 => 32676,
    1095 => 32676,
    1096 => 32677,
    1097 => 32677,
    1098 => 32678,
    1099 => 32678,
    1100 => 32678,
    1101 => 32679,
    1102 => 32679,
    1103 => 32680,
    1104 => 32680,
    1105 => 32681,
    1106 => 32681,
    1107 => 32682,
    1108 => 32682,
    1109 => 32683,
    1110 => 32683,
    1111 => 32684,
    1112 => 32684,
    1113 => 32684,
    1114 => 32685,
    1115 => 32685,
    1116 => 32686,
    1117 => 32686,
    1118 => 32687,
    1119 => 32687,
    1120 => 32687,
    1121 => 32688,
    1122 => 32688,
    1123 => 32689,
    1124 => 32689,
    1125 => 32690,
    1126 => 32690,
    1127 => 32690,
    1128 => 32691,
    1129 => 32691,
    1130 => 32692,
    1131 => 32692,
    1132 => 32692,
    1133 => 32693,
    1134 => 32693,
    1135 => 32694,
    1136 => 32694,
    1137 => 32694,
    1138 => 32695,
    1139 => 32695,
    1140 => 32696,
    1141 => 32696,
    1142 => 32696,
    1143 => 32697,
    1144 => 32697,
    1145 => 32697,
    1146 => 32698,
    1147 => 32698,
    1148 => 32699,
    1149 => 32699,
    1150 => 32699,
    1151 => 32700,
    1152 => 32700,
    1153 => 32700,
    1154 => 32701,
    1155 => 32701,
    1156 => 32701,
    1157 => 32702,
    1158 => 32702,
    1159 => 32702,
    1160 => 32703,
    1161 => 32703,
    1162 => 32704,
    1163 => 32704,
    1164 => 32704,
    1165 => 32705,
    1166 => 32705,
    1167 => 32705,
    1168 => 32706,
    1169 => 32706,
    1170 => 32706,
    1171 => 32706,
    1172 => 32707,
    1173 => 32707,
    1174 => 32707,
    1175 => 32708,
    1176 => 32708,
    1177 => 32708,
    1178 => 32709,
    1179 => 32709,
    1180 => 32709,
    1181 => 32710,
    1182 => 32710,
    1183 => 32710,
    1184 => 32711,
    1185 => 32711,
    1186 => 32711,
    1187 => 32711,
    1188 => 32712,
    1189 => 32712,
    1190 => 32712,
    1191 => 32713,
    1192 => 32713,
    1193 => 32713,
    1194 => 32714,
    1195 => 32714,
    1196 => 32714,
    1197 => 32714,
    1198 => 32715,
    1199 => 32715,
    1200 => 32715,
    1201 => 32715,
    1202 => 32716,
    1203 => 32716,
    1204 => 32716,
    1205 => 32717,
    1206 => 32717,
    1207 => 32717,
    1208 => 32717,
    1209 => 32718,
    1210 => 32718,
    1211 => 32718,
    1212 => 32718,
    1213 => 32719,
    1214 => 32719,
    1215 => 32719,
    1216 => 32719,
    1217 => 32720,
    1218 => 32720,
    1219 => 32720,
    1220 => 32720,
    1221 => 32721,
    1222 => 32721,
    1223 => 32721,
    1224 => 32721,
    1225 => 32722,
    1226 => 32722,
    1227 => 32722,
    1228 => 32722,
    1229 => 32723,
    1230 => 32723,
    1231 => 32723,
    1232 => 32723,
    1233 => 32724,
    1234 => 32724,
    1235 => 32724,
    1236 => 32724,
    1237 => 32725,
    1238 => 32725,
    1239 => 32725,
    1240 => 32725,
    1241 => 32725,
    1242 => 32726,
    1243 => 32726,
    1244 => 32726,
    1245 => 32726,
    1246 => 32727,
    1247 => 32727,
    1248 => 32727,
    1249 => 32727,
    1250 => 32727,
    1251 => 32728,
    1252 => 32728,
    1253 => 32728,
    1254 => 32728,
    1255 => 32728,
    1256 => 32729,
    1257 => 32729,
    1258 => 32729,
    1259 => 32729,
    1260 => 32729,
    1261 => 32730,
    1262 => 32730,
    1263 => 32730,
    1264 => 32730,
    1265 => 32730,
    1266 => 32731,
    1267 => 32731,
    1268 => 32731,
    1269 => 32731,
    1270 => 32731,
    1271 => 32732,
    1272 => 32732,
    1273 => 32732,
    1274 => 32732,
    1275 => 32732,
    1276 => 32733,
    1277 => 32733,
    1278 => 32733,
    1279 => 32733,
    1280 => 32733,
    1281 => 32733,
    1282 => 32734,
    1283 => 32734,
    1284 => 32734,
    1285 => 32734,
    1286 => 32734,
    1287 => 32735,
    1288 => 32735,
    1289 => 32735,
    1290 => 32735,
    1291 => 32735,
    1292 => 32735,
    1293 => 32736,
    1294 => 32736,
    1295 => 32736,
    1296 => 32736,
    1297 => 32736,
    1298 => 32736,
    1299 => 32737,
    1300 => 32737,
    1301 => 32737,
    1302 => 32737,
    1303 => 32737,
    1304 => 32737,
    1305 => 32738,
    1306 => 32738,
    1307 => 32738,
    1308 => 32738,
    1309 => 32738,
    1310 => 32738,
    1311 => 32738,
    1312 => 32739,
    1313 => 32739,
    1314 => 32739,
    1315 => 32739,
    1316 => 32739,
    1317 => 32739,
    1318 => 32740,
    1319 => 32740,
    1320 => 32740,
    1321 => 32740,
    1322 => 32740,
    1323 => 32740,
    1324 => 32740,
    1325 => 32741,
    1326 => 32741,
    1327 => 32741,
    1328 => 32741,
    1329 => 32741,
    1330 => 32741,
    1331 => 32741,
    1332 => 32742,
    1333 => 32742,
    1334 => 32742,
    1335 => 32742,
    1336 => 32742,
    1337 => 32742,
    1338 => 32742,
    1339 => 32742,
    1340 => 32743,
    1341 => 32743,
    1342 => 32743,
    1343 => 32743,
    1344 => 32743,
    1345 => 32743,
    1346 => 32743,
    1347 => 32743,
    1348 => 32744,
    1349 => 32744,
    1350 => 32744,
    1351 => 32744,
    1352 => 32744,
    1353 => 32744,
    1354 => 32744,
    1355 => 32744,
    1356 => 32745,
    1357 => 32745,
    1358 => 32745,
    1359 => 32745,
    1360 => 32745,
    1361 => 32745,
    1362 => 32745,
    1363 => 32745,
    1364 => 32746,
    1365 => 32746,
    1366 => 32746,
    1367 => 32746,
    1368 => 32746,
    1369 => 32746,
    1370 => 32746,
    1371 => 32746,
    1372 => 32746,
    1373 => 32747,
    1374 => 32747,
    1375 => 32747,
    1376 => 32747,
    1377 => 32747,
    1378 => 32747,
    1379 => 32747,
    1380 => 32747,
    1381 => 32747,
    1382 => 32748,
    1383 => 32748,
    1384 => 32748,
    1385 => 32748,
    1386 => 32748,
    1387 => 32748,
    1388 => 32748,
    1389 => 32748,
    1390 => 32748,
    1391 => 32748,
    1392 => 32749,
    1393 => 32749,
    1394 => 32749,
    1395 => 32749,
    1396 => 32749,
    1397 => 32749,
    1398 => 32749,
    1399 => 32749,
    1400 => 32749,
    1401 => 32749,
    1402 => 32749,
    1403 => 32750,
    1404 => 32750,
    1405 => 32750,
    1406 => 32750,
    1407 => 32750,
    1408 => 32750,
    1409 => 32750,
    1410 => 32750,
    1411 => 32750,
    1412 => 32750,
    1413 => 32750,
    1414 => 32751,
    1415 => 32751,
    1416 => 32751,
    1417 => 32751,
    1418 => 32751,
    1419 => 32751,
    1420 => 32751,
    1421 => 32751,
    1422 => 32751,
    1423 => 32751,
    1424 => 32751,
    1425 => 32752,
    1426 => 32752,
    1427 => 32752,
    1428 => 32752,
    1429 => 32752,
    1430 => 32752,
    1431 => 32752,
    1432 => 32752,
    1433 => 32752,
    1434 => 32752,
    1435 => 32752,
    1436 => 32752,
    1437 => 32752,
    1438 => 32753,
    1439 => 32753,
    1440 => 32753,
    1441 => 32753,
    1442 => 32753,
    1443 => 32753,
    1444 => 32753,
    1445 => 32753,
    1446 => 32753,
    1447 => 32753,
    1448 => 32753,
    1449 => 32753,
    1450 => 32753,
    1451 => 32754,
    1452 => 32754,
    1453 => 32754,
    1454 => 32754,
    1455 => 32754,
    1456 => 32754,
    1457 => 32754,
    1458 => 32754,
    1459 => 32754,
    1460 => 32754,
    1461 => 32754,
    1462 => 32754,
    1463 => 32754,
    1464 => 32754,
    1465 => 32755,
    1466 => 32755,
    1467 => 32755,
    1468 => 32755,
    1469 => 32755,
    1470 => 32755,
    1471 => 32755,
    1472 => 32755,
    1473 => 32755,
    1474 => 32755,
    1475 => 32755,
    1476 => 32755,
    1477 => 32755,
    1478 => 32755,
    1479 => 32755,
    1480 => 32755,
    1481 => 32756,
    1482 => 32756,
    1483 => 32756,
    1484 => 32756,
    1485 => 32756,
    1486 => 32756,
    1487 => 32756,
    1488 => 32756,
    1489 => 32756,
    1490 => 32756,
    1491 => 32756,
    1492 => 32756,
    1493 => 32756,
    1494 => 32756,
    1495 => 32756,
    1496 => 32756,
    1497 => 32756,
    1498 => 32757,
    1499 => 32757,
    1500 => 32757,
    1501 => 32757,
    1502 => 32757,
    1503 => 32757,
    1504 => 32757,
    1505 => 32757,
    1506 => 32757,
    1507 => 32757,
    1508 => 32757,
    1509 => 32757,
    1510 => 32757,
    1511 => 32757,
    1512 => 32757,
    1513 => 32757,
    1514 => 32757,
    1515 => 32757,
    1516 => 32758,
    1517 => 32758,
    1518 => 32758,
    1519 => 32758,
    1520 => 32758,
    1521 => 32758,
    1522 => 32758,
    1523 => 32758,
    1524 => 32758,
    1525 => 32758,
    1526 => 32758,
    1527 => 32758,
    1528 => 32758,
    1529 => 32758,
    1530 => 32758,
    1531 => 32758,
    1532 => 32758,
    1533 => 32758,
    1534 => 32758,
    1535 => 32758,
    1536 => 32758,
    1537 => 32759,
    1538 => 32759,
    1539 => 32759,
    1540 => 32759,
    1541 => 32759,
    1542 => 32759,
    1543 => 32759,
    1544 => 32759,
    1545 => 32759,
    1546 => 32759,
    1547 => 32759,
    1548 => 32759,
    1549 => 32759,
    1550 => 32759,
    1551 => 32759,
    1552 => 32759,
    1553 => 32759,
    1554 => 32759,
    1555 => 32759,
    1556 => 32759,
    1557 => 32759,
    1558 => 32759,
    1559 => 32759,
    1560 => 32760,
    1561 => 32760,
    1562 => 32760,
    1563 => 32760,
    1564 => 32760,
    1565 => 32760,
    1566 => 32760,
    1567 => 32760,
    1568 => 32760,
    1569 => 32760,
    1570 => 32760,
    1571 => 32760,
    1572 => 32760,
    1573 => 32760,
    1574 => 32760,
    1575 => 32760,
    1576 => 32760,
    1577 => 32760,
    1578 => 32760,
    1579 => 32760,
    1580 => 32760,
    1581 => 32760,
    1582 => 32760,
    1583 => 32760,
    1584 => 32760,
    1585 => 32760,
    1586 => 32760,
    1587 => 32761,
    1588 => 32761,
    1589 => 32761,
    1590 => 32761,
    1591 => 32761,
    1592 => 32761,
    1593 => 32761,
    1594 => 32761,
    1595 => 32761,
    1596 => 32761,
    1597 => 32761,
    1598 => 32761,
    1599 => 32761,
    1600 => 32761,
    1601 => 32761,
    1602 => 32761,
    1603 => 32761,
    1604 => 32761,
    1605 => 32761,
    1606 => 32761,
    1607 => 32761,
    1608 => 32761,
    1609 => 32761,
    1610 => 32761,
    1611 => 32761,
    1612 => 32761,
    1613 => 32761,
    1614 => 32761,
    1615 => 32761,
    1616 => 32761,
    1617 => 32761,
    1618 => 32762,
    1619 => 32762,
    1620 => 32762,
    1621 => 32762,
    1622 => 32762,
    1623 => 32762,
    1624 => 32762,
    1625 => 32762,
    1626 => 32762,
    1627 => 32762,
    1628 => 32762,
    1629 => 32762,
    1630 => 32762,
    1631 => 32762,
    1632 => 32762,
    1633 => 32762,
    1634 => 32762,
    1635 => 32762,
    1636 => 32762,
    1637 => 32762,
    1638 => 32762,
    1639 => 32762,
    1640 => 32762,
    1641 => 32762,
    1642 => 32762,
    1643 => 32762,
    1644 => 32762,
    1645 => 32762,
    1646 => 32762,
    1647 => 32762,
    1648 => 32762,
    1649 => 32762,
    1650 => 32762,
    1651 => 32762,
    1652 => 32762,
    1653 => 32762,
    1654 => 32762,
    1655 => 32763,
    1656 => 32763,
    1657 => 32763,
    1658 => 32763,
    1659 => 32763,
    1660 => 32763,
    1661 => 32763,
    1662 => 32763,
    1663 => 32763,
    1664 => 32763,
    1665 => 32763,
    1666 => 32763,
    1667 => 32763,
    1668 => 32763,
    1669 => 32763,
    1670 => 32763,
    1671 => 32763,
    1672 => 32763,
    1673 => 32763,
    1674 => 32763,
    1675 => 32763,
    1676 => 32763,
    1677 => 32763,
    1678 => 32763,
    1679 => 32763,
    1680 => 32763,
    1681 => 32763,
    1682 => 32763,
    1683 => 32763,
    1684 => 32763,
    1685 => 32763,
    1686 => 32763,
    1687 => 32763,
    1688 => 32763,
    1689 => 32763,
    1690 => 32763,
    1691 => 32763,
    1692 => 32763,
    1693 => 32763,
    1694 => 32763,
    1695 => 32763,
    1696 => 32763,
    1697 => 32763,
    1698 => 32763,
    1699 => 32763,
    1700 => 32763,
    1701 => 32763,
    1702 => 32764,
    1703 => 32764,
    1704 => 32764,
    1705 => 32764,
    1706 => 32764,
    1707 => 32764,
    1708 => 32764,
    1709 => 32764,
    1710 => 32764,
    1711 => 32764,
    1712 => 32764,
    1713 => 32764,
    1714 => 32764,
    1715 => 32764,
    1716 => 32764,
    1717 => 32764,
    1718 => 32764,
    1719 => 32764,
    1720 => 32764,
    1721 => 32764,
    1722 => 32764,
    1723 => 32764,
    1724 => 32764,
    1725 => 32764,
    1726 => 32764,
    1727 => 32764,
    1728 => 32764,
    1729 => 32764,
    1730 => 32764,
    1731 => 32764,
    1732 => 32764,
    1733 => 32764,
    1734 => 32764,
    1735 => 32764,
    1736 => 32764,
    1737 => 32764,
    1738 => 32764,
    1739 => 32764,
    1740 => 32764,
    1741 => 32764,
    1742 => 32764,
    1743 => 32764,
    1744 => 32764,
    1745 => 32764,
    1746 => 32764,
    1747 => 32764,
    1748 => 32764,
    1749 => 32764,
    1750 => 32764,
    1751 => 32764,
    1752 => 32764,
    1753 => 32764,
    1754 => 32764,
    1755 => 32764,
    1756 => 32764,
    1757 => 32764,
    1758 => 32764,
    1759 => 32764,
    1760 => 32764,
    1761 => 32764,
    1762 => 32764,
    1763 => 32764,
    1764 => 32764,
    1765 => 32765,
    1766 => 32765,
    1767 => 32765,
    1768 => 32765,
    1769 => 32765,
    1770 => 32765,
    1771 => 32765,
    1772 => 32765,
    1773 => 32765,
    1774 => 32765,
    1775 => 32765,
    1776 => 32765,
    1777 => 32765,
    1778 => 32765,
    1779 => 32765,
    1780 => 32765,
    1781 => 32765,
    1782 => 32765,
    1783 => 32765,
    1784 => 32765,
    1785 => 32765,
    1786 => 32765,
    1787 => 32765,
    1788 => 32765,
    1789 => 32765,
    1790 => 32765,
    1791 => 32765,
    1792 => 32765,
    1793 => 32765,
    1794 => 32765,
    1795 => 32765,
    1796 => 32765,
    1797 => 32765,
    1798 => 32765,
    1799 => 32765,
    1800 => 32765,
    1801 => 32765,
    1802 => 32765,
    1803 => 32765,
    1804 => 32765,
    1805 => 32765,
    1806 => 32765,
    1807 => 32765,
    1808 => 32765,
    1809 => 32765,
    1810 => 32765,
    1811 => 32765,
    1812 => 32765,
    1813 => 32765,
    1814 => 32765,
    1815 => 32765,
    1816 => 32765,
    1817 => 32765,
    1818 => 32765,
    1819 => 32765,
    1820 => 32765,
    1821 => 32765,
    1822 => 32765,
    1823 => 32765,
    1824 => 32765,
    1825 => 32765,
    1826 => 32765,
    1827 => 32765,
    1828 => 32765,
    1829 => 32765,
    1830 => 32765,
    1831 => 32765,
    1832 => 32765,
    1833 => 32765,
    1834 => 32765,
    1835 => 32765,
    1836 => 32765,
    1837 => 32765,
    1838 => 32765,
    1839 => 32765,
    1840 => 32765,
    1841 => 32765,
    1842 => 32765,
    1843 => 32765,
    1844 => 32765,
    1845 => 32765,
    1846 => 32765,
    1847 => 32765,
    1848 => 32765,
    1849 => 32765,
    1850 => 32765,
    1851 => 32765,
    1852 => 32765,
    1853 => 32765,
    1854 => 32765,
    1855 => 32765,
    1856 => 32765,
    1857 => 32765,
    1858 => 32765,
    1859 => 32765,
    1860 => 32766,
    1861 => 32766,
    1862 => 32766,
    1863 => 32766,
    1864 => 32766,
    1865 => 32766,
    1866 => 32766,
    1867 => 32766,
    1868 => 32766,
    1869 => 32766,
    1870 => 32766,
    1871 => 32766,
    1872 => 32766,
    1873 => 32766,
    1874 => 32766,
    1875 => 32766,
    1876 => 32766,
    1877 => 32766,
    1878 => 32766,
    1879 => 32766,
    1880 => 32766,
    1881 => 32766,
    1882 => 32766,
    1883 => 32766,
    1884 => 32766,
    1885 => 32766,
    1886 => 32766,
    1887 => 32766,
    1888 => 32766,
    1889 => 32766,
    1890 => 32766,
    1891 => 32766,
    1892 => 32766,
    1893 => 32766,
    1894 => 32766,
    1895 => 32766,
    1896 => 32766,
    1897 => 32766,
    1898 => 32766,
    1899 => 32766,
    1900 => 32766,
    1901 => 32766,
    1902 => 32766,
    1903 => 32766,
    1904 => 32766,
    1905 => 32766,
    1906 => 32766,
    1907 => 32766,
    1908 => 32766,
    1909 => 32766,
    1910 => 32766,
    1911 => 32766,
    1912 => 32766,
    1913 => 32766,
    1914 => 32766,
    1915 => 32766,
    1916 => 32766,
    1917 => 32766,
    1918 => 32766,
    1919 => 32766,
    1920 => 32766,
    1921 => 32766,
    1922 => 32766,
    1923 => 32766,
    1924 => 32766,
    1925 => 32766,
    1926 => 32766,
    1927 => 32766,
    1928 => 32766,
    1929 => 32766,
    1930 => 32766,
    1931 => 32766,
    1932 => 32766,
    1933 => 32766,
    1934 => 32766,
    1935 => 32766,
    1936 => 32766,
    1937 => 32766,
    1938 => 32766,
    1939 => 32766,
    1940 => 32766,
    1941 => 32766,
    1942 => 32766,
    1943 => 32766,
    1944 => 32766,
    1945 => 32766,
    1946 => 32766,
    1947 => 32766,
    1948 => 32766,
    1949 => 32766,
    1950 => 32766,
    1951 => 32766,
    1952 => 32766,
    1953 => 32766,
    1954 => 32766,
    1955 => 32766,
    1956 => 32766,
    1957 => 32766,
    1958 => 32766,
    1959 => 32766,
    1960 => 32766,
    1961 => 32766,
    1962 => 32766,
    1963 => 32766,
    1964 => 32766,
    1965 => 32766,
    1966 => 32766,
    1967 => 32766,
    1968 => 32766,
    1969 => 32766,
    1970 => 32766,
    1971 => 32766,
    1972 => 32766,
    1973 => 32766,
    1974 => 32766,
    1975 => 32766,
    1976 => 32766,
    1977 => 32766,
    1978 => 32766,
    1979 => 32766,
    1980 => 32766,
    1981 => 32766,
    1982 => 32766,
    1983 => 32766,
    1984 => 32766,
    1985 => 32766,
    1986 => 32766,
    1987 => 32766,
    1988 => 32766,
    1989 => 32766,
    1990 => 32766,
    1991 => 32766,
    1992 => 32766,
    1993 => 32766,
    1994 => 32766,
    1995 => 32766,
    1996 => 32766,
    1997 => 32766,
    1998 => 32766,
    1999 => 32766,
    2000 => 32766,
    2001 => 32766,
    2002 => 32766,
    2003 => 32766,
    2004 => 32766,
    2005 => 32766,
    2006 => 32766,
    2007 => 32766,
    2008 => 32766,
    2009 => 32766,
    2010 => 32766,
    2011 => 32766,
    2012 => 32766,
    2013 => 32766,
    2014 => 32766,
    2015 => 32766,
    2016 => 32766,
    2017 => 32766,
    2018 => 32766,
    2019 => 32766,
    2020 => 32766,
    2021 => 32766,
    2022 => 32766,
    2023 => 32766,
    2024 => 32766,
    2025 => 32766,
    2026 => 32766,
    2027 => 32766,
    2028 => 32766,
    2029 => 32766,
    2030 => 32766,
    2031 => 32766,
    2032 => 32766,
    2033 => 32766,
    2034 => 32766,
    2035 => 32766,
    2036 => 32766,
    2037 => 32766,
    2038 => 32766,
    2039 => 32766,
    2040 => 32766,
    2041 => 32766,
    2042 => 32766,
    2043 => 32766,
    2044 => 32766,
    2045 => 32766,
    2046 => 32766,
    2047 => 32766
);

begin
  dds_out <= std_logic_vector(TO_SIGNED(LUT(TO_INTEGER(unsigned(address))),16));
end rtl;
